`include "FPA.v"

module top;
	
	reg [31:0] a,b;
	wire [31:0] sum;
	
	initial
		begin
			$dumpfile("FPA_32bit.vcd");
			$dumpvars(0,top);
		end
	
	initial
		begin
			//A = 9.75, B = 0.5625
			a = 32'b01000001000111000000000000000000;
			b = 32'b00111111000100000000000000000000;
			
			//A = 0, B = 0.5625
			#100
			a = 32'b00000000000000000000000000000000;
			b = 32'b00111111000100000000000000000000;
			
			//A = 9.75, B = Infinity
			#100
			a = 32'b01000001000111000000000000000000;
			b = 32'b01111111100000000000000000000000;
			
			//A = 9.75, B = -9.75
			#100
			a = 32'b01000001000111000000000000000000;
			b = 32'b11000001000111000000000000000000;
			
		end
	
	FPA_32BIT fp_adder(a,b,sum);
	
	initial
		$monitor("\n\t\tX1 = %b\n\t\tX2 = %b\n\n\t\tX3 = %b\n" ,a,b,sum);
	
endmodule
