module parallelprefix(
	input x0_j_1,
	input x1_j_1,
	input x0_j,
	input x1_j,
	output reg y0,
	output reg y1
	);
	
	always @(x0_j_1,x1_j_1,x0_j,x1_j)
		begin
			if((x0_j_1^x1_j_1)==1'b0)
				begin
					assign y0=x0_j_1;
					assign y1=x1_j_1;
				end
			else
				begin
					assign y0=x0_j;
					assign y1=x1_j;
				end
		end

endmodule

module recursive_doubling(
	input [63:0] x0,
	input [63:0] x1,
	output [63:0] f0,
	output [63:0] f1
	);
	
	wire [63:0] y0,y1;
	wire [63:0] z0,z1;
	wire [63:0] p0,p1;
	wire [63:0] q0,q1;
	wire [63:0] r0,r1;
	
	parallelprefix kpg0(x0[63],x1[63],x0[62],x1[62],y0[63],y1[63]);
	parallelprefix kpg1(x0[62],x1[62],x0[61],x1[61],y0[62],y1[62]);
	parallelprefix kpg2(x0[61],x1[61],x0[60],x1[60],y0[61],y1[61]);
	parallelprefix kpg3(x0[60],x1[60],x0[59],x1[59],y0[60],y1[60]);
	parallelprefix kpg4(x0[59],x1[59],x0[58],x1[58],y0[59],y1[59]);
	parallelprefix kpg5(x0[58],x1[58],x0[57],x1[57],y0[58],y1[58]);
	parallelprefix kpg6(x0[57],x1[57],x0[56],x1[56],y0[57],y1[57]);
	parallelprefix kpg7(x0[56],x1[56],x0[55],x1[55],y0[56],y1[56]);
	parallelprefix kpg8(x0[55],x1[55],x0[54],x1[54],y0[55],y1[55]);
	parallelprefix kpg9(x0[54],x1[54],x0[53],x1[53],y0[54],y1[54]);
	parallelprefix kpg10(x0[53],x1[53],x0[52],x1[52],y0[53],y1[53]);
	parallelprefix kpg11(x0[52],x1[52],x0[51],x1[51],y0[52],y1[52]);
	parallelprefix kpg12(x0[51],x1[51],x0[50],x1[50],y0[51],y1[51]);
	parallelprefix kpg13(x0[50],x1[50],x0[49],x1[49],y0[50],y1[50]);
	parallelprefix kpg14(x0[49],x1[49],x0[48],x1[48],y0[49],y1[49]);
	parallelprefix kpg15(x0[48],x1[48],x0[47],x1[47],y0[48],y1[48]);
	parallelprefix kpg16(x0[47],x1[47],x0[46],x1[46],y0[47],y1[47]);
	parallelprefix kpg17(x0[46],x1[46],x0[45],x1[45],y0[46],y1[46]);
	parallelprefix kpg18(x0[45],x1[45],x0[44],x1[44],y0[45],y1[45]);
	parallelprefix kpg19(x0[44],x1[44],x0[43],x1[43],y0[44],y1[44]);
	parallelprefix kpg20(x0[43],x1[43],x0[42],x1[42],y0[43],y1[43]);
	parallelprefix kpg21(x0[42],x1[42],x0[41],x1[41],y0[42],y1[42]);
	parallelprefix kpg22(x0[41],x1[41],x0[40],x1[40],y0[41],y1[41]);
	parallelprefix kpg23(x0[40],x1[40],x0[39],x1[39],y0[40],y1[40]);
	parallelprefix kpg24(x0[39],x1[39],x0[38],x1[38],y0[39],y1[39]);
	parallelprefix kpg25(x0[38],x1[38],x0[37],x1[37],y0[38],y1[38]);
	parallelprefix kpg26(x0[37],x1[37],x0[36],x1[36],y0[37],y1[37]);
	parallelprefix kpg27(x0[36],x1[36],x0[35],x1[35],y0[36],y1[36]);
	parallelprefix kpg28(x0[35],x1[35],x0[34],x1[34],y0[35],y1[35]);
	parallelprefix kpg29(x0[34],x1[34],x0[33],x1[33],y0[34],y1[34]);
	parallelprefix kpg30(x0[33],x1[33],x0[32],x1[32],y0[33],y1[33]);
	parallelprefix kpg31(x0[32],x1[32],x0[31],x1[31],y0[32],y1[32]);
	parallelprefix kpg32(x0[31],x1[31],x0[30],x1[30],y0[31],y1[31]);
	parallelprefix kpg33(x0[30],x1[30],x0[29],x1[29],y0[30],y1[30]);
	parallelprefix kpg34(x0[29],x1[29],x0[28],x1[28],y0[29],y1[29]);
	parallelprefix kpg35(x0[28],x1[28],x0[27],x1[27],y0[28],y1[28]);
	parallelprefix kpg36(x0[27],x1[27],x0[26],x1[26],y0[27],y1[27]);
	parallelprefix kpg37(x0[26],x1[26],x0[25],x1[25],y0[26],y1[26]);
	parallelprefix kpg38(x0[25],x1[25],x0[24],x1[24],y0[25],y1[25]);
	parallelprefix kpg39(x0[24],x1[24],x0[23],x1[23],y0[24],y1[24]);
	parallelprefix kpg40(x0[23],x1[23],x0[22],x1[22],y0[23],y1[23]);
	parallelprefix kpg41(x0[22],x1[22],x0[21],x1[21],y0[22],y1[22]);
	parallelprefix kpg42(x0[21],x1[21],x0[20],x1[20],y0[21],y1[21]);
	parallelprefix kpg43(x0[20],x1[20],x0[19],x1[19],y0[20],y1[20]);
	parallelprefix kpg44(x0[19],x1[19],x0[18],x1[18],y0[19],y1[19]);
	parallelprefix kpg45(x0[18],x1[18],x0[17],x1[17],y0[18],y1[18]);
	parallelprefix kpg46(x0[17],x1[17],x0[16],x1[16],y0[17],y1[17]);
	parallelprefix kpg47(x0[16],x1[16],x0[15],x1[15],y0[16],y1[16]);
	parallelprefix kpg48(x0[15],x1[15],x0[14],x1[14],y0[15],y1[15]);
	parallelprefix kpg49(x0[14],x1[14],x0[13],x1[13],y0[14],y1[14]);
	parallelprefix kpg50(x0[13],x1[13],x0[12],x1[12],y0[13],y1[13]);
	parallelprefix kpg51(x0[12],x1[12],x0[11],x1[11],y0[12],y1[12]);
	parallelprefix kpg52(x0[11],x1[11],x0[10],x1[10],y0[11],y1[11]);
	parallelprefix kpg53(x0[10],x1[10],x0[9],x1[9],y0[10],y1[10]);
	parallelprefix kpg54(x0[9],x1[9],x0[8],x1[8],y0[9],y1[9]);
	parallelprefix kpg55(x0[8],x1[8],x0[7],x1[7],y0[8],y1[8]);
	parallelprefix kpg56(x0[7],x1[7],x0[6],x1[6],y0[7],y1[7]);
	parallelprefix kpg57(x0[6],x1[6],x0[5],x1[5],y0[6],y1[6]);
	parallelprefix kpg58(x0[5],x1[5],x0[4],x1[4],y0[5],y1[5]);
	parallelprefix kpg59(x0[4],x1[4],x0[3],x1[3],y0[4],y1[4]);
	parallelprefix kpg60(x0[3],x1[3],x0[2],x1[2],y0[3],y1[3]);
	parallelprefix kpg61(x0[2],x1[2],x0[1],x1[1],y0[2],y1[2]);
	parallelprefix kpg62(x0[1],x1[1],x0[0],x1[0],y0[1],y1[1]);
	parallelprefix kpg63(x0[0],x1[0],1'b0,1'b0,y0[0],y1[0]);
	
	
	parallelprefix kpg64(y0[63],y1[63],y0[61],y1[61],z0[63],z1[63]);
	parallelprefix kpg65(y0[62],y1[62],y0[60],y1[60],z0[62],z1[62]);
	parallelprefix kpg66(y0[61],y1[61],y0[59],y1[59],z0[61],z1[61]);
	parallelprefix kpg67(y0[60],y1[60],y0[58],y1[58],z0[60],z1[60]);
	parallelprefix kpg68(y0[59],y1[59],y0[57],y1[57],z0[59],z1[59]);
	parallelprefix kpg69(y0[58],y1[58],y0[56],y1[56],z0[58],z1[58]);
	parallelprefix kpg70(y0[57],y1[57],y0[55],y1[55],z0[57],z1[57]);
	parallelprefix kpg71(y0[56],y1[56],y0[54],y1[54],z0[56],z1[56]);
	parallelprefix kpg72(y0[55],y1[55],y0[53],y1[53],z0[55],z1[55]);
	parallelprefix kpg73(y0[54],y1[54],y0[52],y1[52],z0[54],z1[54]);
	parallelprefix kpg74(y0[53],y1[53],y0[51],y1[51],z0[53],z1[53]);
	parallelprefix kpg75(y0[52],y1[52],y0[50],y1[50],z0[52],z1[52]);
	parallelprefix kpg76(y0[51],y1[51],y0[49],y1[49],z0[51],z1[51]);
	parallelprefix kpg77(y0[50],y1[50],y0[48],y1[48],z0[50],z1[50]);
	parallelprefix kpg78(y0[49],y1[49],y0[47],y1[47],z0[49],z1[49]);
	parallelprefix kpg79(y0[48],y1[48],y0[46],y1[46],z0[48],z1[48]);
	parallelprefix kpg80(y0[47],y1[47],y0[45],y1[45],z0[47],z1[47]);
	parallelprefix kpg81(y0[46],y1[46],y0[44],y1[44],z0[46],z1[46]);
	parallelprefix kpg82(y0[45],y1[45],y0[43],y1[43],z0[45],z1[45]);
	parallelprefix kpg83(y0[44],y1[44],y0[42],y1[42],z0[44],z1[44]);
	parallelprefix kpg84(y0[43],y1[43],y0[41],y1[41],z0[43],z1[43]);
	parallelprefix kpg85(y0[42],y1[42],y0[40],y1[40],z0[42],z1[42]);
	parallelprefix kpg86(y0[41],y1[41],y0[39],y1[39],z0[41],z1[41]);
	parallelprefix kpg87(y0[40],y1[40],y0[38],y1[38],z0[40],z1[40]);
	parallelprefix kpg88(y0[39],y1[39],y0[37],y1[37],z0[39],z1[39]);
	parallelprefix kpg89(y0[38],y1[38],y0[36],y1[36],z0[38],z1[38]);
	parallelprefix kpg90(y0[37],y1[37],y0[35],y1[35],z0[37],z1[37]);
	parallelprefix kpg91(y0[36],y1[36],y0[34],y1[34],z0[36],z1[36]);
	parallelprefix kpg92(y0[35],y1[35],y0[33],y1[33],z0[35],z1[35]);
	parallelprefix kpg93(y0[34],y1[34],y0[32],y1[32],z0[34],z1[34]);
	parallelprefix kpg94(y0[33],y1[33],y0[31],y1[31],z0[33],z1[33]);
	parallelprefix kpg95(y0[32],y1[32],y0[30],y1[30],z0[32],z1[32]);
	parallelprefix kpg96(y0[31],y1[31],y0[29],y1[29],z0[31],z1[31]);
	parallelprefix kpg97(y0[30],y1[30],y0[28],y1[28],z0[30],z1[30]);
	parallelprefix kpg98(y0[29],y1[29],y0[27],y1[27],z0[29],z1[29]);
	parallelprefix kpg99(y0[28],y1[28],y0[26],y1[26],z0[28],z1[28]);
	parallelprefix kpg100(y0[27],y1[27],y0[25],y1[25],z0[27],z1[27]);
	parallelprefix kpg101(y0[26],y1[26],y0[24],y1[24],z0[26],z1[26]);
	parallelprefix kpg102(y0[25],y1[25],y0[23],y1[23],z0[25],z1[25]);
	parallelprefix kpg103(y0[24],y1[24],y0[22],y1[22],z0[24],z1[24]);
	parallelprefix kpg104(y0[23],y1[23],y0[21],y1[21],z0[23],z1[23]);
	parallelprefix kpg105(y0[22],y1[22],y0[20],y1[20],z0[22],z1[22]);
	parallelprefix kpg106(y0[21],y1[21],y0[19],y1[19],z0[21],z1[21]);
	parallelprefix kpg107(y0[20],y1[20],y0[18],y1[18],z0[20],z1[20]);
	parallelprefix kpg108(y0[19],y1[19],y0[17],y1[17],z0[19],z1[19]);
	parallelprefix kpg109(y0[18],y1[18],y0[16],y1[16],z0[18],z1[18]);
	parallelprefix kpg110(y0[17],y1[17],y0[15],y1[15],z0[17],z1[17]);
	parallelprefix kpg111(y0[16],y1[16],y0[14],y1[14],z0[16],z1[16]);
	parallelprefix kpg112(y0[15],y1[15],y0[13],y1[13],z0[15],z1[15]);
	parallelprefix kpg113(y0[14],y1[14],y0[12],y1[12],z0[14],z1[14]);
	parallelprefix kpg114(y0[13],y1[13],y0[11],y1[11],z0[13],z1[13]);
	parallelprefix kpg115(y0[12],y1[12],y0[10],y1[10],z0[12],z1[12]);
	parallelprefix kpg116(y0[11],y1[11],y0[9],y1[9],z0[11],z1[11]);
	parallelprefix kpg117(y0[10],y1[10],y0[8],y1[8],z0[10],z1[10]);
	parallelprefix kpg118(y0[9],y1[9],y0[7],y1[7],z0[9],z1[9]);
	parallelprefix kpg119(y0[8],y1[8],y0[6],y1[6],z0[8],z1[8]);
	parallelprefix kpg120(y0[7],y1[7],y0[5],y1[5],z0[7],z1[7]);
	parallelprefix kpg121(y0[6],y1[6],y0[4],y1[4],z0[6],z1[6]);
	parallelprefix kpg122(y0[5],y1[5],y0[3],y1[3],z0[5],z1[5]);
	parallelprefix kpg123(y0[4],y1[4],y0[2],y1[2],z0[4],z1[4]);
	parallelprefix kpg124(y0[3],y1[3],y0[1],y1[1],z0[3],z1[3]);
	parallelprefix kpg125(y0[2],y1[2],y0[0],y1[0],z0[2],z1[2]);
	parallelprefix kpg126(y0[1],y1[1],1'b0,1'b0,z0[1],z1[1]);
	parallelprefix kpg127(y0[0],y1[0],y0[0],y1[0],z0[0],z1[0]);
	
	
	parallelprefix kpg_0(z0[63],z1[63],z0[59],z1[59],p0[63],p1[63]);
	parallelprefix kpg_1(z0[62],z1[62],z0[58],z1[58],p0[62],p1[62]);
	parallelprefix kpg_2(z0[61],z1[61],z0[57],z1[57],p0[61],p1[61]);
	parallelprefix kpg_3(z0[60],z1[60],z0[56],z1[56],p0[60],p1[60]);
	parallelprefix kpg_4(z0[59],z1[59],z0[55],z1[55],p0[59],p1[59]);
	parallelprefix kpg_5(z0[58],z1[58],z0[54],z1[54],p0[58],p1[58]);
	parallelprefix kpg_6(z0[57],z1[57],z0[53],z1[53],p0[57],p1[57]);
	parallelprefix kpg_7(z0[56],z1[56],z0[52],z1[52],p0[56],p1[56]);
	parallelprefix kpg_8(z0[55],z1[55],z0[51],z1[51],p0[55],p1[55]);
	parallelprefix kpg_9(z0[54],z1[54],z0[50],z1[50],p0[54],p1[54]);
	parallelprefix kpg_10(z0[53],z1[53],z0[49],z1[49],p0[53],p1[53]);
	parallelprefix kpg_11(z0[52],z1[52],z0[48],z1[48],p0[52],p1[52]);
	parallelprefix kpg_12(z0[51],z1[51],z0[47],z1[47],p0[51],p1[51]);
	parallelprefix kpg_13(z0[50],z1[50],z0[46],z1[46],p0[50],p1[50]);
	parallelprefix kpg_14(z0[49],z1[49],z0[45],z1[45],p0[49],p1[49]);
	parallelprefix kpg_15(z0[48],z1[48],z0[44],z1[44],p0[48],p1[48]);
	parallelprefix kpg_16(z0[47],z1[47],z0[43],z1[43],p0[47],p1[47]);
	parallelprefix kpg_17(z0[46],z1[46],z0[42],z1[42],p0[46],p1[46]);
	parallelprefix kpg_18(z0[45],z1[45],z0[41],z1[41],p0[45],p1[45]);
	parallelprefix kpg_19(z0[44],z1[44],z0[40],z1[40],p0[44],p1[44]);
	parallelprefix kpg_20(z0[43],z1[43],z0[39],z1[39],p0[43],p1[43]);
	parallelprefix kpg_21(z0[42],z1[42],z0[38],z1[38],p0[42],p1[42]);
	parallelprefix kpg_22(z0[41],z1[41],z0[37],z1[37],p0[41],p1[41]);
	parallelprefix kpg_23(z0[40],z1[40],z0[36],z1[36],p0[40],p1[40]);
	parallelprefix kpg_24(z0[39],z1[39],z0[35],z1[35],p0[39],p1[39]);
	parallelprefix kpg_25(z0[38],z1[38],z0[34],z1[34],p0[38],p1[38]);
	parallelprefix kpg_26(z0[37],z1[37],z0[33],z1[33],p0[37],p1[37]);
	parallelprefix kpg_27(z0[36],z1[36],z0[32],z1[32],p0[36],p1[36]);
	parallelprefix kpg_28(z0[35],z1[35],z0[31],z1[31],p0[35],p1[35]);
	parallelprefix kpg_29(z0[34],z1[34],z0[30],z1[30],p0[34],p1[34]);
	parallelprefix kpg_30(z0[33],z1[33],z0[29],z1[29],p0[33],p1[33]);
	parallelprefix kpg_31(z0[32],z1[32],z0[28],z1[28],p0[32],p1[32]);
	parallelprefix kpg_32(z0[31],z1[31],z0[27],z1[27],p0[31],p1[31]);
	parallelprefix kpg_33(z0[30],z1[30],z0[26],z1[26],p0[30],p1[30]);
	parallelprefix kpg_34(z0[29],z1[29],z0[25],z1[25],p0[29],p1[29]);
	parallelprefix kpg_35(z0[28],z1[28],z0[24],z1[24],p0[28],p1[28]);
	parallelprefix kpg_36(z0[27],z1[27],z0[23],z1[23],p0[27],p1[27]);
	parallelprefix kpg_37(z0[26],z1[26],z0[22],z1[22],p0[26],p1[26]);
	parallelprefix kpg_38(z0[25],z1[25],z0[21],z1[21],p0[25],p1[25]);
	parallelprefix kpg_39(z0[24],z1[24],z0[20],z1[20],p0[24],p1[24]);
	parallelprefix kpg_40(z0[23],z1[23],z0[19],z1[19],p0[23],p1[23]);
	parallelprefix kpg_41(z0[22],z1[22],z0[18],z1[18],p0[22],p1[22]);
	parallelprefix kpg_42(z0[21],z1[21],z0[17],z1[17],p0[21],p1[21]);
	parallelprefix kpg_43(z0[20],z1[20],z0[16],z1[16],p0[20],p1[20]);
	parallelprefix kpg_44(z0[19],z1[19],z0[15],z1[15],p0[19],p1[19]);
	parallelprefix kpg_45(z0[18],z1[18],z0[14],z1[14],p0[18],p1[18]);
	parallelprefix kpg_46(z0[17],z1[17],z0[13],z1[13],p0[17],p1[17]);
	parallelprefix kpg_47(z0[16],z1[16],z0[12],z1[12],p0[16],p1[16]);
	parallelprefix kpg_48(z0[15],z1[15],z0[11],z1[11],p0[15],p1[15]);
	parallelprefix kpg_49(z0[14],z1[14],z0[10],z1[10],p0[14],p1[14]);
	parallelprefix kpg_50(z0[13],z1[13],z0[9],z1[9],p0[13],p1[13]);
	parallelprefix kpg_51(z0[12],z1[12],z0[8],z1[8],p0[12],p1[12]);
	parallelprefix kpg_52(z0[11],z1[11],z0[7],z1[7],p0[11],p1[11]);
	parallelprefix kpg_53(z0[10],z1[10],z0[6],z1[6],p0[10],p1[10]);
	parallelprefix kpg_54(z0[9],z1[9],z0[5],z1[5],p0[9],p1[9]);
	parallelprefix kpg_55(z0[8],z1[8],z0[4],z1[4],p0[8],p1[8]);
	parallelprefix kpg_56(z0[7],z1[7],z0[3],z1[3],p0[7],p1[7]);
	parallelprefix kpg_57(z0[6],z1[6],z0[2],z1[2],p0[6],p1[6]);
	parallelprefix kpg_58(z0[5],z1[5],z0[1],z1[1],p0[5],p1[5]);
	parallelprefix kpg_59(z0[4],z1[4],z0[0],z1[0],p0[4],p1[4]);
	parallelprefix kpg_60(z0[3],z1[3],1'b0,1'b0,p0[3],p1[3]);
	parallelprefix kpg_61(z0[2],z1[2],z0[2],z1[2],p0[2],p1[2]);
	parallelprefix kpg_62(z0[1],z1[1],z0[1],z1[1],p0[1],p1[1]);
	parallelprefix kpg_63(z0[0],z1[0],z0[0],z1[0],p0[0],p1[0]);

	
	parallelprefix kpg_64(p0[63],p1[63],p0[55],p1[55],q0[63],q1[63]);
	parallelprefix kpg_65(p0[62],p1[62],p0[54],p1[54],q0[62],q1[62]);
	parallelprefix kpg_66(p0[61],p1[61],p0[53],p1[53],q0[61],q1[61]);
	parallelprefix kpg_67(p0[60],p1[60],p0[52],p1[52],q0[60],q1[60]);
	parallelprefix kpg_68(p0[59],p1[59],p0[51],p1[51],q0[59],q1[59]);
	parallelprefix kpg_69(p0[58],p1[58],p0[50],p1[50],q0[58],q1[58]);
	parallelprefix kpg_70(p0[57],p1[57],p0[49],p1[49],q0[57],q1[57]);
	parallelprefix kpg_71(p0[56],p1[56],p0[48],p1[48],q0[56],q1[56]);
	parallelprefix kpg_72(p0[55],p1[55],p0[47],p1[47],q0[55],q1[55]);
	parallelprefix kpg_73(p0[54],p1[54],p0[46],p1[46],q0[54],q1[54]);
	parallelprefix kpg_74(p0[53],p1[53],p0[45],p1[45],q0[53],q1[53]);
	parallelprefix kpg_75(p0[52],p1[52],p0[44],p1[44],q0[52],q1[52]);
	parallelprefix kpg_76(p0[51],p1[51],p0[43],p1[43],q0[51],q1[51]);
	parallelprefix kpg_77(p0[50],p1[50],p0[42],p1[42],q0[50],q1[50]);
	parallelprefix kpg_78(p0[49],p1[49],p0[41],p1[41],q0[49],q1[49]);
	parallelprefix kpg_79(p0[48],p1[48],p0[40],p1[40],q0[48],q1[48]);
	parallelprefix kpg_80(p0[47],p1[47],p0[39],p1[39],q0[47],q1[47]);
	parallelprefix kpg_81(p0[46],p1[46],p0[38],p1[38],q0[46],q1[46]);
	parallelprefix kpg_82(p0[45],p1[45],p0[37],p1[37],q0[45],q1[45]);
	parallelprefix kpg_83(p0[44],p1[44],p0[36],p1[36],q0[44],q1[44]);
	parallelprefix kpg_84(p0[43],p1[43],p0[35],p1[35],q0[43],q1[43]);
	parallelprefix kpg_85(p0[42],p1[42],p0[34],p1[34],q0[42],q1[42]);
	parallelprefix kpg_86(p0[41],p1[41],p0[33],p1[33],q0[41],q1[41]);
	parallelprefix kpg_87(p0[40],p1[40],p0[32],p1[32],q0[40],q1[40]);
	parallelprefix kpg_88(p0[39],p1[39],p0[31],p1[31],q0[39],q1[39]);
	parallelprefix kpg_89(p0[38],p1[38],p0[30],p1[30],q0[38],q1[38]);
	parallelprefix kpg_90(p0[37],p1[37],p0[29],p1[29],q0[37],q1[37]);
	parallelprefix kpg_91(p0[36],p1[36],p0[28],p1[28],q0[36],q1[36]);
	parallelprefix kpg_92(p0[35],p1[35],p0[27],p1[27],q0[35],q1[35]);
	parallelprefix kpg_93(p0[34],p1[34],p0[26],p1[26],q0[34],q1[34]);
	parallelprefix kpg_94(p0[33],p1[33],p0[25],p1[25],q0[33],q1[33]);
	parallelprefix kpg_95(p0[32],p1[32],p0[24],p1[24],q0[32],q1[32]);
	parallelprefix kpg_96(p0[31],p1[31],p0[23],p1[23],q0[31],q1[31]);
	parallelprefix kpg_97(p0[30],p1[30],p0[22],p1[22],q0[30],q1[30]);
	parallelprefix kpg_98(p0[29],p1[29],p0[21],p1[21],q0[29],q1[29]);
	parallelprefix kpg_99(p0[28],p1[28],p0[20],p1[20],q0[28],q1[28]);
	parallelprefix kpg_100(p0[27],p1[27],p0[19],p1[19],q0[27],q1[27]);
	parallelprefix kpg_101(p0[26],p1[26],p0[18],p1[18],q0[26],q1[26]);
	parallelprefix kpg_102(p0[25],p1[25],p0[17],p1[17],q0[25],q1[25]);
	parallelprefix kpg_103(p0[24],p1[24],p0[18],p1[16],q0[24],q1[24]);
	parallelprefix kpg_104(p0[23],p1[23],p0[15],p1[15],q0[23],q1[23]);
	parallelprefix kpg_105(p0[22],p1[22],p0[14],p1[14],q0[22],q1[22]);
	parallelprefix kpg_106(p0[21],p1[21],p0[13],p1[13],q0[21],q1[21]);
	parallelprefix kpg_107(p0[20],p1[20],p0[12],p1[12],q0[20],q1[20]);
	parallelprefix kpg_108(p0[19],p1[19],p0[11],p1[11],q0[29],q1[19]);
	parallelprefix kpg_109(p0[18],p1[18],p0[10],p1[10],q0[18],q1[18]);
	parallelprefix kpg_110(p0[17],p1[17],p0[9],p1[9],q0[17],q1[17]);
	parallelprefix kpg_111(p0[16],p1[16],p0[8],p1[8],q0[16],q1[16]);
	parallelprefix kpg_112(p0[15],p1[15],p0[7],p1[7],q0[15],q1[15]);
	parallelprefix kpg_113(p0[14],p1[14],p0[6],p1[6],q0[14],q1[14]);
	parallelprefix kpg_114(p0[13],p1[13],p0[5],p1[5],q0[13],q1[13]);
	parallelprefix kpg_115(p0[12],p1[12],p0[4],p1[4],q0[12],q1[12]);
	parallelprefix kpg_116(p0[11],p1[11],p0[3],p1[3],q0[11],q1[11]);
	parallelprefix kpg_117(p0[10],p1[10],p0[2],p1[2],q0[10],q1[10]);
	parallelprefix kpg_118(p0[9],p1[9],p0[1],p1[1],q0[9],q1[9]);
	parallelprefix kpg_119(p0[8],p1[8],p0[0],p1[0],q0[8],q1[8]);
	parallelprefix kpg_120(p0[7],p1[7],1'b0,1'b0,q0[7],q1[7]);
	parallelprefix kpg_121(p0[6],p1[6],p0[6],p1[6],q0[6],q1[6]);
	parallelprefix kpg_122(p0[5],p1[5],p0[5],p1[5],q0[5],q1[5]);
	parallelprefix kpg_123(p0[4],p1[4],p0[4],p1[4],q0[4],q1[4]);
	parallelprefix kpg_124(p0[3],p1[3],p0[3],p1[3],q0[3],q1[3]);
	parallelprefix kpg_125(p0[2],p1[2],p0[2],p1[2],q0[2],q1[2]);
	parallelprefix kpg_126(p0[1],p1[1],p0[1],p1[1],q0[1],q1[1]);
	parallelprefix kpg_127(p0[0],p1[0],p0[0],p1[0],q0[0],q1[0]);


	parallelprefix kpg_00(q0[63],q1[63],q0[47],q1[47],r0[63],r1[63]);
	parallelprefix kpg_01(q0[62],q1[62],q0[46],q1[46],r0[62],r1[62]);
	parallelprefix kpg_02(q0[61],q1[61],q0[45],q1[45],r0[61],r1[61]);
	parallelprefix kpg_03(q0[60],q1[60],q0[44],q1[44],r0[60],r1[60]);
	parallelprefix kpg_04(q0[59],q1[59],q0[43],q1[43],r0[59],r1[59]);
	parallelprefix kpg_05(q0[58],q1[58],q0[42],q1[42],r0[58],r1[58]);
	parallelprefix kpg_06(q0[57],q1[57],q0[41],q1[41],r0[57],r1[57]);
	parallelprefix kpg_07(q0[56],q1[56],q0[40],q1[40],r0[56],r1[56]);
	parallelprefix kpg_08(q0[55],q1[55],q0[39],q1[39],r0[55],r1[55]);
	parallelprefix kpg_09(q0[54],q1[54],q0[38],q1[38],r0[54],r1[54]);
	parallelprefix kpg_010(q0[53],q1[53],q0[37],q1[37],r0[53],r1[53]);
	parallelprefix kpg_011(q0[52],q1[52],q0[36],q1[36],r0[52],r1[52]);
	parallelprefix kpg_012(q0[51],q1[51],q0[35],q1[35],r0[51],r1[51]);
	parallelprefix kpg_013(q0[50],q1[50],q0[34],q1[34],r0[50],r1[50]);
	parallelprefix kpg_014(q0[49],q1[49],q0[33],q1[33],r0[49],r1[49]);
	parallelprefix kpg_015(q0[48],q1[48],q0[32],q1[32],r0[48],r1[48]);
	parallelprefix kpg_016(q0[47],q1[47],q0[31],q1[31],r0[47],r1[47]);
	parallelprefix kpg_017(q0[46],q1[46],q0[30],q1[30],r0[46],r1[46]);
	parallelprefix kpg_018(q0[45],q1[45],q0[29],q1[29],r0[45],r1[45]);
	parallelprefix kpg_019(q0[44],q1[44],q0[28],q1[28],r0[44],r1[44]);
	parallelprefix kpg_020(q0[43],q1[43],q0[27],q1[27],r0[43],r1[43]);
	parallelprefix kpg_021(q0[42],q1[42],q0[26],q1[26],r0[42],r1[42]);
	parallelprefix kpg_022(q0[41],q1[41],q0[25],q1[25],r0[41],r1[41]);
	parallelprefix kpg_023(q0[40],q1[40],q0[24],q1[24],r0[40],r1[40]);
	parallelprefix kpg_024(q0[39],q1[39],q0[23],q1[23],r0[39],r1[39]);
	parallelprefix kpg_025(q0[38],q1[38],q0[22],q1[22],r0[38],r1[38]);
	parallelprefix kpg_026(q0[37],q1[37],q0[21],q1[21],r0[37],r1[37]);
	parallelprefix kpg_027(q0[36],q1[36],q0[20],q1[20],r0[36],r1[36]);
	parallelprefix kpg_028(q0[35],q1[35],q0[19],q1[19],r0[35],r1[35]);
	parallelprefix kpg_029(q0[34],q1[34],q0[18],q1[18],r0[34],r1[34]);
	parallelprefix kpg_030(q0[33],q1[33],q0[17],q1[17],r0[33],r1[33]);
	parallelprefix kpg_031(q0[32],q1[32],q0[16],q1[16],r0[32],r1[32]);
	parallelprefix kpg_032(q0[31],q1[31],q0[15],q1[15],r0[31],r1[31]);
	parallelprefix kpg_033(q0[30],q1[30],q0[14],q1[14],r0[30],r1[30]);
	parallelprefix kpg_034(q0[29],q1[29],q0[13],q1[13],r0[29],r1[29]);
	parallelprefix kpg_035(q0[28],q1[28],q0[12],q1[12],r0[28],r1[28]);
	parallelprefix kpg_036(q0[27],q1[27],q0[11],q1[11],r0[27],r1[27]);
	parallelprefix kpg_037(q0[26],q1[26],q0[10],q1[10],r0[26],r1[26]);
	parallelprefix kpg_038(q0[25],q1[25],q0[9],q1[9],r0[25],r1[25]);
	parallelprefix kpg_039(q0[24],q1[24],q0[8],q1[8],r0[24],r1[24]);
	parallelprefix kpg_040(q0[23],q1[23],q0[7],q1[7],r0[23],r1[23]);
	parallelprefix kpg_041(q0[22],q1[22],q0[6],q1[6],r0[22],r1[22]);
	parallelprefix kpg_042(q0[21],q1[21],q0[5],q1[5],r0[21],r1[21]);
	parallelprefix kpg_043(q0[20],q1[20],q0[4],q1[4],r0[20],r1[20]);
	parallelprefix kpg_044(q0[19],q1[19],q0[3],q1[3],r0[19],r1[19]);
	parallelprefix kpg_045(q0[18],q1[18],q0[2],q1[2],r0[18],r1[18]);
	parallelprefix kpg_046(q0[17],q1[17],q0[1],q1[1],r0[17],r1[17]);
	parallelprefix kpg_047(q0[16],q1[16],q0[0],q1[0],r0[16],r1[16]);
	parallelprefix kpg_048(q0[15],q1[15],1'b0,1'b0,r0[15],r1[15]);
	parallelprefix kpg_049(q0[14],q1[14],q0[14],q1[14],r0[14],r1[14]);
	parallelprefix kpg_050(q0[13],q1[13],q0[13],q1[13],r0[13],r1[13]);
	parallelprefix kpg_051(q0[12],q1[12],q0[12],q1[12],r0[12],r1[12]);
	parallelprefix kpg_052(q0[11],q1[11],q0[11],q1[11],r0[11],r1[11]);
	parallelprefix kpg_053(q0[10],q1[10],q0[10],q1[10],r0[10],r1[10]);
	parallelprefix kpg_054(q0[9],q1[9],q0[9],q1[9],r0[9],r1[9]);
	parallelprefix kpg_055(q0[8],q1[8],q0[8],q1[8],r0[8],r1[8]);
	parallelprefix kpg_056(q0[7],q1[7],q0[7],q1[7],r0[7],r1[7]);
	parallelprefix kpg_057(q0[6],q1[6],q0[6],q1[6],r0[6],r1[6]);
	parallelprefix kpg_058(q0[5],q1[5],q0[5],q1[5],r0[5],r1[5]);
	parallelprefix kpg_059(q0[4],q1[4],q0[4],q1[4],r0[4],r1[4]);
	parallelprefix kpg_060(q0[3],q1[3],q0[3],q1[3],r0[3],r1[3]);
	parallelprefix kpg_061(q0[2],q1[2],q0[2],q1[2],r0[2],r1[2]);
	parallelprefix kpg_062(q0[1],q1[1],q0[1],q1[1],r0[1],r1[1]);
	parallelprefix kpg_063(q0[0],q1[0],q0[0],q1[0],r0[0],r1[0]);


	parallelprefix kpg_064(r0[63],r1[63],r0[31],r1[31],f0[63],f1[63]);
	parallelprefix kpg_065(r0[62],r1[62],r0[30],r1[30],f0[62],f1[62]);
	parallelprefix kpg_066(r0[61],r1[61],r0[29],r1[29],f0[61],f1[61]);
	parallelprefix kpg_067(r0[60],r1[60],r0[28],r1[28],f0[60],f1[60]);
	parallelprefix kpg_068(r0[59],r1[59],r0[27],r1[27],f0[59],f1[59]);
	parallelprefix kpg_069(r0[58],r1[58],r0[26],r1[26],f0[58],f1[58]);
	parallelprefix kpg_070(r0[57],r1[57],r0[25],r1[25],f0[57],f1[57]);
	parallelprefix kpg_071(r0[56],r1[56],r0[24],r1[24],f0[56],f1[56]);
	parallelprefix kpg_072(r0[55],r1[55],r0[23],r1[23],f0[55],f1[55]);
	parallelprefix kpg_073(r0[54],r1[54],r0[22],r1[22],f0[54],f1[54]);
	parallelprefix kpg_074(r0[53],r1[53],r0[21],r1[21],f0[53],f1[53]);
	parallelprefix kpg_075(r0[52],r1[52],r0[20],r1[20],f0[52],f1[52]);
	parallelprefix kpg_076(r0[51],r1[51],r0[19],r1[19],f0[51],f1[51]);
	parallelprefix kpg_077(r0[50],r1[50],r0[18],r1[18],f0[50],f1[50]);
	parallelprefix kpg_078(r0[49],r1[49],r0[17],r1[17],f0[49],f1[49]);
	parallelprefix kpg_079(r0[48],r1[48],r0[16],r1[16],f0[48],f1[48]);
	parallelprefix kpg_080(r0[47],r1[47],r0[15],r1[15],f0[47],f1[47]);
	parallelprefix kpg_081(r0[46],r1[46],r0[14],r1[14],f0[46],f1[46]);
	parallelprefix kpg_082(r0[45],r1[45],r0[13],r1[13],f0[45],f1[45]);
	parallelprefix kpg_083(r0[44],r1[44],r0[12],r1[12],f0[44],f1[44]);
	parallelprefix kpg_084(r0[43],r1[43],r0[11],r1[11],f0[43],f1[43]);
	parallelprefix kpg_085(r0[42],r1[42],r0[10],r1[10],f0[42],f1[42]);
	parallelprefix kpg_086(r0[41],r1[41],r0[9],r1[9],f0[41],f1[41]);
	parallelprefix kpg_087(r0[40],r1[40],r0[8],r1[8],f0[40],f1[40]);
	parallelprefix kpg_088(r0[39],r1[39],r0[7],r1[7],f0[39],f1[39]);
	parallelprefix kpg_089(r0[38],r1[38],r0[6],r1[6],f0[38],f1[38]);
	parallelprefix kpg_090(r0[37],r1[37],r0[5],r1[5],f0[37],f1[37]);
	parallelprefix kpg_091(r0[36],r1[36],r0[4],r1[4],f0[36],f1[36]);
	parallelprefix kpg_092(r0[35],r1[35],r0[3],r1[3],f0[35],f1[35]);
	parallelprefix kpg_093(r0[34],r1[34],r0[2],r1[2],f0[34],f1[34]);
	parallelprefix kpg_094(r0[33],r1[33],r0[1],r1[1],f0[33],f1[33]);
	parallelprefix kpg_095(r0[32],r1[32],r0[0],r1[0],f0[32],f1[32]);
	parallelprefix kpg_096(r0[31],r1[31],1'b0,1'b0,f0[31],f1[31]);
	parallelprefix kpg_097(r0[30],r1[30],r0[30],r1[30],f0[30],f1[30]);
	parallelprefix kpg_098(r0[29],r1[29],r0[29],r1[29],f0[29],f1[29]);
	parallelprefix kpg_099(r0[28],r1[28],r0[28],r1[28],f0[28],f1[28]);
	parallelprefix kpg_0100(r0[27],r1[27],r0[27],r1[27],f0[27],f1[27]);
	parallelprefix kpg_0101(r0[26],r1[26],r0[26],r1[26],f0[26],f1[26]);
	parallelprefix kpg_0102(r0[25],r1[25],r0[25],r1[25],f0[25],f1[25]);
	parallelprefix kpg_0103(r0[24],r1[24],r0[24],r1[24],f0[24],f1[24]);
	parallelprefix kpg_0104(r0[23],r1[23],r0[23],r1[23],f0[23],f1[23]);
	parallelprefix kpg_0105(r0[22],r1[22],r0[22],r1[22],f0[22],f1[22]);
	parallelprefix kpg_0106(r0[21],r1[21],r0[21],r1[21],f0[21],f1[21]);
	parallelprefix kpg_0107(r0[20],r1[20],r0[20],r1[20],f0[20],f1[20]);
	parallelprefix kpg_0108(r0[19],r1[19],r0[19],r1[19],f0[19],f1[19]);
	parallelprefix kpg_0109(r0[18],r1[18],r0[18],r1[18],f0[18],f1[18]);
	parallelprefix kpg_0110(r0[17],r1[17],r0[17],r1[17],f0[17],f1[17]);
	parallelprefix kpg_0111(r0[16],r1[16],r0[16],r1[16],f0[16],f1[16]);
	parallelprefix kpg_0112(r0[15],r1[15],r0[15],r1[15],f0[15],f1[15]);
	parallelprefix kpg_0113(r0[14],r1[14],r0[14],r1[14],f0[14],f1[14]);
	parallelprefix kpg_0114(r0[13],r1[13],r0[13],r1[13],f0[13],f1[13]);
	parallelprefix kpg_0115(r0[12],r1[12],r0[12],r1[12],f0[12],f1[12]);
	parallelprefix kpg_0116(r0[11],r1[11],r0[11],r1[11],f0[11],f1[11]);
	parallelprefix kpg_0117(r0[10],r1[10],r0[10],r1[10],f0[10],f1[10]);
	parallelprefix kpg_0118(r0[9],r1[9],r0[9],r1[9],f0[9],f1[9]);
	parallelprefix kpg_0119(r0[8],r1[8],r0[8],r1[8],f0[8],f1[8]);
	parallelprefix kpg_0120(r0[7],r1[7],r0[7],r1[7],f0[7],f1[7]);
	parallelprefix kpg_0121(r0[6],r1[6],r0[6],r1[6],f0[6],f1[6]);
	parallelprefix kpg_0122(r0[5],r1[5],r0[5],r1[5],f0[5],f1[5]);
	parallelprefix kpg_0123(r0[4],r1[4],r0[4],r1[4],f0[4],f1[4]);
	parallelprefix kpg_0124(r0[3],r1[3],r0[3],r1[3],f0[3],f1[3]);
	parallelprefix kpg_0125(r0[2],r1[2],r0[2],r1[2],f0[2],f1[2]);
	parallelprefix kpg_0126(r0[1],r1[1],r0[1],r1[1],f0[1],f1[1]);
	parallelprefix kpg_0127(r0[0],r1[0],r0[0],r1[0],f0[0],f1[0]);


endmodule

module Adder_64bit(
	input [63:0] a,
	input [63:0] b,
	output [63:0] sum
	);
	
	wire [63:0] sum_without_carry,carry;
	wire [63:0] x0,x1;
	wire [63:0] f0,f1;
	
	assign sum_without_carry[0]=a[0]^b[0];
	assign sum_without_carry[1]=a[1]^b[1];
	assign sum_without_carry[2]=a[2]^b[2];
	assign sum_without_carry[3]=a[3]^b[3];
	assign sum_without_carry[4]=a[4]^b[4];
	assign sum_without_carry[5]=a[5]^b[5];
	assign sum_without_carry[6]=a[6]^b[6];
	assign sum_without_carry[7]=a[7]^b[7];
	assign sum_without_carry[8]=a[8]^b[8];
	assign sum_without_carry[9]=a[9]^b[9];
	assign sum_without_carry[10]=a[10]^b[10];
	assign sum_without_carry[11]=a[11]^b[11];
	assign sum_without_carry[12]=a[12]^b[12];
	assign sum_without_carry[13]=a[13]^b[13];
	assign sum_without_carry[14]=a[14]^b[14];
	assign sum_without_carry[15]=a[15]^b[15];
	assign sum_without_carry[16]=a[16]^b[16];
	assign sum_without_carry[17]=a[17]^b[17];
	assign sum_without_carry[18]=a[18]^b[18];
	assign sum_without_carry[19]=a[19]^b[19];
	assign sum_without_carry[20]=a[20]^b[20];
	assign sum_without_carry[21]=a[21]^b[21];
	assign sum_without_carry[22]=a[22]^b[22];
	assign sum_without_carry[23]=a[23]^b[23];
	assign sum_without_carry[24]=a[24]^b[24];
	assign sum_without_carry[25]=a[25]^b[25];
	assign sum_without_carry[26]=a[26]^b[26];
	assign sum_without_carry[27]=a[27]^b[27];
	assign sum_without_carry[28]=a[28]^b[28];
	assign sum_without_carry[29]=a[29]^b[29];
	assign sum_without_carry[30]=a[30]^b[30];
	assign sum_without_carry[31]=a[31]^b[31];
	assign sum_without_carry[32]=a[32]^b[32];
	assign sum_without_carry[33]=a[33]^b[33];
	assign sum_without_carry[34]=a[34]^b[34];
	assign sum_without_carry[35]=a[35]^b[35];
	assign sum_without_carry[36]=a[36]^b[36];
	assign sum_without_carry[37]=a[37]^b[37];
	assign sum_without_carry[38]=a[38]^b[38];
	assign sum_without_carry[39]=a[39]^b[39];
	assign sum_without_carry[40]=a[40]^b[40];
	assign sum_without_carry[41]=a[41]^b[41];
	assign sum_without_carry[42]=a[42]^b[42];
	assign sum_without_carry[43]=a[43]^b[43];
	assign sum_without_carry[44]=a[44]^b[44];
	assign sum_without_carry[45]=a[45]^b[45];
	assign sum_without_carry[46]=a[46]^b[46];
	assign sum_without_carry[47]=a[47]^b[47];
	assign sum_without_carry[48]=a[48]^b[48];
	assign sum_without_carry[49]=a[49]^b[49];
	assign sum_without_carry[50]=a[50]^b[50];
	assign sum_without_carry[51]=a[51]^b[51];
	assign sum_without_carry[52]=a[52]^b[52];
	assign sum_without_carry[53]=a[53]^b[53];
	assign sum_without_carry[54]=a[54]^b[54];
	assign sum_without_carry[55]=a[55]^b[55];
	assign sum_without_carry[56]=a[56]^b[56];
	assign sum_without_carry[57]=a[57]^b[57];
	assign sum_without_carry[58]=a[58]^b[58];
	assign sum_without_carry[59]=a[59]^b[59];
	assign sum_without_carry[60]=a[60]^b[60];
	assign sum_without_carry[61]=a[61]^b[61];
	assign sum_without_carry[62]=a[62]^b[62];
	assign sum_without_carry[63]=a[63]^b[63];
	
	
	assign x0[0]=a[0]|b[0];
	assign x1[0]=a[0]&b[0];
	assign x0[1]=a[1]|b[1];
	assign x1[1]=a[1]&b[1];
	assign x0[2]=a[2]|b[2];
	assign x1[2]=a[2]&b[2];
	assign x0[3]=a[3]|b[3];
	assign x1[3]=a[3]&b[3];
	assign x0[4]=a[4]|b[4];
	assign x1[4]=a[4]&b[4];
	assign x0[5]=a[5]|b[5];
	assign x1[5]=a[5]&b[5];
	assign x0[6]=a[6]|b[6];
	assign x1[6]=a[6]&b[6];
	assign x0[7]=a[7]|b[7];
	assign x1[7]=a[7]&b[7];
	assign x0[8]=a[8]|b[8];
	assign x1[8]=a[8]&b[8];
	assign x0[9]=a[9]|b[9];
	assign x1[9]=a[9]&b[9];
	assign x0[10]=a[10]|b[10];
	assign x1[10]=a[10]&b[10];
	assign x0[11]=a[11]|b[11];
	assign x1[11]=a[11]&b[11];
	assign x0[12]=a[12]|b[12];
	assign x1[12]=a[12]&b[12];
	assign x0[13]=a[13]|b[13];
	assign x1[13]=a[13]&b[13];
	assign x0[14]=a[14]|b[14];
	assign x1[14]=a[14]&b[14];
	assign x0[15]=a[15]|b[15];
	assign x1[15]=a[15]&b[15];
	assign x0[16]=a[16]|b[16];
	assign x1[16]=a[16]&b[16];
	assign x0[17]=a[17]|b[17];
	assign x1[17]=a[17]&b[17];
	assign x0[18]=a[18]|b[18];
	assign x1[18]=a[18]&b[18];
	assign x0[19]=a[19]|b[19];
	assign x1[19]=a[19]&b[19];
	assign x0[20]=a[20]|b[20];
	assign x1[20]=a[20]&b[20];
	assign x0[21]=a[21]|b[21];
	assign x1[21]=a[21]&b[21];
	assign x0[22]=a[22]|b[22];
	assign x1[22]=a[22]&b[22];
	assign x0[23]=a[23]|b[23];
	assign x1[23]=a[23]&b[23];
	assign x0[24]=a[24]|b[24];
	assign x1[24]=a[24]&b[24];
	assign x0[25]=a[25]|b[25];
	assign x1[25]=a[25]&b[25];
	assign x0[26]=a[26]|b[26];
	assign x1[26]=a[26]&b[26];
	assign x1[27]=a[27]&b[27];
	assign x0[27]=a[27]|b[27];
	assign x0[28]=a[28]|b[28];
	assign x1[28]=a[28]&b[28];
	assign x1[29]=a[29]&b[29];
	assign x0[29]=a[29]|b[29];
	assign x0[30]=a[30]|b[30];
	assign x1[30]=a[30]&b[30];
	assign x0[31]=a[31]|b[31];
	assign x1[31]=a[31]&b[31];
	assign x0[32]=a[32]|b[32];
	assign x1[32]=a[32]&b[32];
	assign x0[33]=a[33]|b[33];
	assign x1[33]=a[33]&b[33];
	assign x0[34]=a[34]|b[34];
	assign x1[34]=a[34]&b[34];
	assign x0[35]=a[35]|b[35];
	assign x1[35]=a[35]&b[35];
	assign x0[36]=a[36]|b[36];
	assign x1[36]=a[36]&b[36];
	assign x0[37]=a[37]|b[37];
	assign x1[37]=a[37]&b[37];
	assign x0[38]=a[38]|b[38];
	assign x1[38]=a[38]&b[38];
	assign x0[39]=a[39]|b[39];
	assign x1[39]=a[39]&b[39];
	assign x0[40]=a[40]|b[40];
	assign x1[40]=a[40]&b[40];
	assign x0[41]=a[41]|b[41];
	assign x1[41]=a[41]&b[41];
	assign x0[42]=a[42]|b[42];
	assign x1[42]=a[42]&b[42];
	assign x0[43]=a[43]|b[43];
	assign x1[43]=a[43]&b[43];
	assign x0[44]=a[44]|b[44];
	assign x1[44]=a[44]&b[44];
	assign x0[45]=a[45]|b[45];
	assign x1[45]=a[45]&b[45];
	assign x0[46]=a[46]|b[46];
	assign x1[46]=a[46]&b[46];
	assign x0[47]=a[47]|b[47];
	assign x1[47]=a[47]&b[47];
	assign x0[48]=a[48]|b[48];
	assign x1[48]=a[48]&b[48];
	assign x0[49]=a[49]|b[49];
	assign x1[49]=a[49]&b[49];
	assign x0[50]=a[50]|b[50];
	assign x1[50]=a[50]&b[50];
	assign x0[51]=a[51]|b[51];
	assign x1[51]=a[51]&b[51];
	assign x0[52]=a[52]|b[52];
	assign x1[52]=a[52]&b[52];
	assign x0[53]=a[53]|b[53];
	assign x1[53]=a[53]&b[53];
	assign x0[54]=a[54]|b[54];
	assign x1[54]=a[54]&b[54];
	assign x0[55]=a[55]|b[55];
	assign x1[55]=a[55]&b[55];
	assign x0[56]=a[56]|b[56];
	assign x1[56]=a[56]&b[56];
	assign x0[57]=a[57]|b[57];
	assign x1[57]=a[57]&b[57];
	assign x0[58]=a[58]|b[58];
	assign x1[58]=a[58]&b[58];
	assign x0[59]=a[59]|b[59];
	assign x1[59]=a[59]&b[59];
	assign x0[60]=a[60]|b[60];
	assign x1[60]=a[60]&b[60];
	assign x0[61]=a[61]|b[61];
	assign x1[61]=a[61]&b[61];
	assign x0[62]=a[62]|b[62];
	assign x1[62]=a[62]&b[62];
	assign x0[63]=a[63]|b[63];
	assign x1[63]=a[63]&b[63];
	
	
	recursive_doubling rd1(x0[63:0],x1[63:0],f0[63:0],f1[63:0]);
	
	assign carry[0]=f1[0]&f0[0];
	assign carry[1]=f1[1]&f0[1];
	assign carry[2]=f1[2]&f0[2];
	assign carry[3]=f1[3]&f0[3];
	assign carry[4]=f1[4]&f0[4];
	assign carry[5]=f1[5]&f0[5];
	assign carry[6]=f1[6]&f0[6];
	assign carry[7]=f1[7]&f0[7];
	assign carry[8]=f1[8]&f0[8];
	assign carry[9]=f1[9]&f0[9];
	assign carry[10]=f1[10]&f0[10];
	assign carry[11]=f1[11]&f0[11];
	assign carry[12]=f1[12]&f0[12];
	assign carry[13]=f1[13]&f0[13];
	assign carry[14]=f1[14]&f0[14];
	assign carry[15]=f1[15]&f0[15];
	assign carry[16]=f1[16]&f0[16];
	assign carry[17]=f1[17]&f0[17];
	assign carry[18]=f1[18]&f0[18];
	assign carry[19]=f1[19]&f0[19];
	assign carry[20]=f1[20]&f0[20];
	assign carry[21]=f1[21]&f0[21];
	assign carry[22]=f1[22]&f0[22];
	assign carry[23]=f1[23]&f0[23];
	assign carry[24]=f1[24]&f0[24];
	assign carry[25]=f1[25]&f0[25];
	assign carry[26]=f1[26]&f0[26];
	assign carry[27]=f1[27]&f0[27];
	assign carry[28]=f1[28]&f0[28];
	assign carry[29]=f1[29]&f0[29];
	assign carry[30]=f1[30]&f0[30];
	assign carry[31]=f1[31]&f0[31];
	assign carry[32]=f1[32]&f0[32];
	assign carry[33]=f1[33]&f0[33];
	assign carry[34]=f1[34]&f0[34];
	assign carry[35]=f1[35]&f0[35];
	assign carry[36]=f1[36]&f0[36];
	assign carry[37]=f1[37]&f0[37];
	assign carry[38]=f1[38]&f0[38];
	assign carry[39]=f1[39]&f0[39];
	assign carry[40]=f1[40]&f0[40];
	assign carry[41]=f1[41]&f0[41];
	assign carry[42]=f1[42]&f0[42];
	assign carry[43]=f1[43]&f0[43];
	assign carry[44]=f1[44]&f0[44];
	assign carry[45]=f1[45]&f0[45];
	assign carry[46]=f1[46]&f0[46];
	assign carry[47]=f1[47]&f0[47];
	assign carry[48]=f1[48]&f0[48];
	assign carry[49]=f1[49]&f0[49];
	assign carry[50]=f1[50]&f0[50];
	assign carry[51]=f1[51]&f0[51];
	assign carry[52]=f1[52]&f0[52];
	assign carry[53]=f1[53]&f0[53];
	assign carry[54]=f1[54]&f0[54];
	assign carry[55]=f1[55]&f0[55];
	assign carry[56]=f1[56]&f0[56];
	assign carry[57]=f1[57]&f0[57];
	assign carry[58]=f1[58]&f0[58];
	assign carry[59]=f1[59]&f0[59];
	assign carry[60]=f1[60]&f0[60];
	assign carry[61]=f1[61]&f0[61];
	assign carry[62]=f1[62]&f0[62];
	assign carry[63]=f1[63]&f0[63];
	
	
	assign sum[0]=sum_without_carry[0];
	assign sum[1]=sum_without_carry[1]^carry[0];
	assign sum[2]=sum_without_carry[2]^carry[1];
	assign sum[3]=sum_without_carry[3]^carry[2];
	assign sum[4]=sum_without_carry[4]^carry[3];
	assign sum[5]=sum_without_carry[5]^carry[4];
	assign sum[6]=sum_without_carry[6]^carry[5];
	assign sum[7]=sum_without_carry[7]^carry[6];
	assign sum[8]=sum_without_carry[8]^carry[7];
	assign sum[9]=sum_without_carry[9]^carry[8];
	assign sum[10]=sum_without_carry[10]^carry[9];
	assign sum[11]=sum_without_carry[11]^carry[10];
	assign sum[12]=sum_without_carry[12]^carry[11];
	assign sum[13]=sum_without_carry[13]^carry[12];
	assign sum[14]=sum_without_carry[14]^carry[13];
	assign sum[15]=sum_without_carry[15]^carry[14];
	assign sum[16]=sum_without_carry[16]^carry[15];
	assign sum[17]=sum_without_carry[17]^carry[16];
	assign sum[18]=sum_without_carry[18]^carry[17];
	assign sum[19]=sum_without_carry[19]^carry[18];
	assign sum[20]=sum_without_carry[20]^carry[19];
	assign sum[21]=sum_without_carry[21]^carry[20];
	assign sum[22]=sum_without_carry[22]^carry[21];
	assign sum[23]=sum_without_carry[23]^carry[22];
	assign sum[24]=sum_without_carry[24]^carry[23];
	assign sum[25]=sum_without_carry[25]^carry[24];
	assign sum[26]=sum_without_carry[26]^carry[25];
	assign sum[27]=sum_without_carry[27]^carry[26];
	assign sum[28]=sum_without_carry[28]^carry[27];
	assign sum[29]=sum_without_carry[29]^carry[28];
	assign sum[30]=sum_without_carry[30]^carry[29];
	assign sum[31]=sum_without_carry[31]^carry[30];
	assign sum[32]=sum_without_carry[32]^carry[31];
	assign sum[33]=sum_without_carry[33]^carry[32];
	assign sum[34]=sum_without_carry[34]^carry[33];
	assign sum[35]=sum_without_carry[35]^carry[34];
	assign sum[36]=sum_without_carry[36]^carry[35];
	assign sum[37]=sum_without_carry[37]^carry[36];
	assign sum[38]=sum_without_carry[38]^carry[37];
	assign sum[39]=sum_without_carry[39]^carry[38];
	assign sum[40]=sum_without_carry[40]^carry[39];
	assign sum[41]=sum_without_carry[41]^carry[40];
	assign sum[42]=sum_without_carry[42]^carry[41];
	assign sum[43]=sum_without_carry[43]^carry[42];
	assign sum[44]=sum_without_carry[44]^carry[43];
	assign sum[45]=sum_without_carry[45]^carry[44];
	assign sum[46]=sum_without_carry[46]^carry[45];
	assign sum[47]=sum_without_carry[47]^carry[46];
	assign sum[48]=sum_without_carry[48]^carry[47];
	assign sum[49]=sum_without_carry[49]^carry[48];
	assign sum[50]=sum_without_carry[50]^carry[49];
	assign sum[51]=sum_without_carry[51]^carry[50];
	assign sum[52]=sum_without_carry[52]^carry[51];
	assign sum[53]=sum_without_carry[53]^carry[52];
	assign sum[54]=sum_without_carry[54]^carry[53];
	assign sum[55]=sum_without_carry[55]^carry[54];
	assign sum[56]=sum_without_carry[56]^carry[55];
	assign sum[57]=sum_without_carry[57]^carry[56];
	assign sum[58]=sum_without_carry[58]^carry[57];
	assign sum[59]=sum_without_carry[59]^carry[58];
	assign sum[60]=sum_without_carry[60]^carry[59];
	assign sum[61]=sum_without_carry[61]^carry[60];
	assign sum[62]=sum_without_carry[62]^carry[61];
	assign sum[63]=sum_without_carry[63]^carry[62];
	
endmodule
