`include "Logic_Unit.v"

module top;
	
	reg [31:0] in1,in2;
    	reg [2:0] select;
	wire [31:0] out;
	
	initial
		begin
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b000;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b001;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b010;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b011;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b100;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b101;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b110;
			
			#10
			in1 = 32'b00000000001000001000111000000000;
			in2 = 32'b00000000000111111000100000000000;
			select = 3'b111;
		end
	
	logic_unit LU(in1,in2,select,out);

	initial
		$monitor("\n\tA = %b\tB = %b\tSelect = %b\tOutput = %b",in1,in2,select,out);
	
endmodule
